module Top (
	input        i_clk,
	input        i_rst,
	input        i_start,
	output [3:0] o_random_out
);

// please check out the working example in lab1 README first

endmodule
