module Rsa256Core (
	input          i_clk,
	input          i_rst,
	input          i_start,
	input  [255:0] i_a,
	input  [255:0] i_e,
	input  [255:0] i_n,
	output [255:0] o_a_pow_e,
	output         o_finished
);

// operations for RSA256 decryption
// namely, the Montgomery algorithm

endmodule
